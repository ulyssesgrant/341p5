// Write a tester here using the readData and writeData tasks

module test
  (output logic clk, rst_L);
  
  
    

endmodule
